module df(q, d, clk, reset);
  output reg q;
  input d, clk, reset;
  always @ (posedge clk or negedge reset)
    begin
      if(~reset) q <= 0;
      else q <= d;
    end
endmodule